module test1(i1,i2,a1);
endmodule
